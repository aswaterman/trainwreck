../vector/vuVXU-Opcode.vh