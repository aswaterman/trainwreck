//**************************************************************************
// Generic Verilog Library: Decoders
//--------------------------------------------------------------------------
// $Id: vcDecoders.v,v 1.1.1.1 2006/02/17 23:57:17 cbatten Exp $
//

//--------------------------------------------------------------------------
// Decoder
//--------------------------------------------------------------------------

module vcDecoder
#(
  parameter W_IN  = 3, 
  parameter W_OUT = 8
) 
(
  input      [W_IN-1:0]  in, 
  output reg [W_OUT-1:0] out
);   

   always @(*) 
   begin
     out     = {W_OUT{1'b0}};
     out[in] = 1'b1;
   end

endmodule
