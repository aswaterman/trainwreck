`ifndef ASIC
`define ASIC
`define CHIP_SMALL

// Define this to disable post-tapeout bug fixes
//`define ST_TAPEOUT_0

`endif
