
module estNormDistP53PosSum108( a, b, out );

    input  [107:0] a, b;
    output [7:0]   out;

    wire [107:0] key;

    assign key = ( a ^ b ) ^ ( ( a | b )<<1 );
    assign out =
          key[107] ?  53
        : key[106] ?  54
        : key[105] ?  55
        : key[104] ?  56
        : key[103] ?  57
        : key[102] ?  58
        : key[101] ?  59
        : key[100] ?  60
        : key[99]  ?  61
        : key[98]  ?  62
        : key[97]  ?  63
        : key[96]  ?  64
        : key[95]  ?  65
        : key[94]  ?  66
        : key[93]  ?  67
        : key[92]  ?  68
        : key[91]  ?  69
        : key[90]  ?  70
        : key[89]  ?  71
        : key[88]  ?  72
        : key[87]  ?  73
        : key[86]  ?  74
        : key[85]  ?  75
        : key[84]  ?  76
        : key[83]  ?  77
        : key[82]  ?  78
        : key[81]  ?  79
        : key[80]  ?  80
        : key[79]  ?  81
        : key[78]  ?  82
        : key[77]  ?  83
        : key[76]  ?  84
        : key[75]  ?  85
        : key[74]  ?  86
        : key[73]  ?  87
        : key[72]  ?  88
        : key[71]  ?  89
        : key[70]  ?  90
        : key[69]  ?  91
        : key[68]  ?  92
        : key[67]  ?  93
        : key[66]  ?  94
        : key[65]  ?  95
        : key[64]  ?  96
        : key[63]  ?  97
        : key[62]  ?  98
        : key[61]  ?  99
        : key[60]  ? 100
        : key[59]  ? 101
        : key[58]  ? 102
        : key[57]  ? 103
        : key[56]  ? 104
        : key[55]  ? 105
        : key[54]  ? 106
        : key[53]  ? 107
        : key[52]  ? 108
        : key[51]  ? 109
        : key[50]  ? 110
        : key[49]  ? 111
        : key[48]  ? 112
        : key[47]  ? 113
        : key[46]  ? 114
        : key[45]  ? 115
        : key[44]  ? 116
        : key[43]  ? 117
        : key[42]  ? 118
        : key[41]  ? 119
        : key[40]  ? 120
        : key[39]  ? 121
        : key[38]  ? 122
        : key[37]  ? 123
        : key[36]  ? 124
        : key[35]  ? 125
        : key[34]  ? 126
        : key[33]  ? 127
        : key[32]  ? 128
        : key[31]  ? 129
        : key[30]  ? 130
        : key[29]  ? 131
        : key[28]  ? 132
        : key[27]  ? 133
        : key[26]  ? 134
        : key[25]  ? 135
        : key[24]  ? 136
        : key[23]  ? 137
        : key[22]  ? 138
        : key[21]  ? 139
        : key[20]  ? 140
        : key[19]  ? 141
        : key[18]  ? 142
        : key[17]  ? 143
        : key[16]  ? 144
        : key[15]  ? 145
        : key[14]  ? 146
        : key[13]  ? 147
        : key[12]  ? 148
        : key[11]  ? 149
        : key[10]  ? 150
        : key[9]   ? 151
        : key[8]   ? 152
        : key[7]   ? 153
        : key[6]   ? 154
        : key[5]   ? 155
        : key[4]   ? 156
        : key[3]   ? 157
        : key[2]   ? 158
        : key[1]   ? 159
        : 160;

endmodule

