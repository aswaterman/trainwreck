../vector/vuVXU-B8-Config.vh